class Test_v3 extends component;
    typedef registry #(Test_v3, "Test_v3") type_id;
endclass // Test_v3
