class TestBad extends component;
    typedef registry #(TestBad, "TestBad") type_id;
endclass // TestBad
