class TestGood extends component;
    typedef registry #(TestGood, "TestGood") type_id;
endclass // TestGood
